.title KiCad schematic
.include "models/C2012X7R2A223K125AE_p.mod"
.include "models/C3216X5R0J107M160AB_p.mod"
.include "models/C3216X7R1H105K160AE_p.mod"
.include "models/C3225X5R1H106K250AB_p.mod"
.include "models/LMZ12003_TRANS.LIB"
XU1 /IN /RON /EN 0 /SS /FB /OUT LMZ12003_TRANS
XU6 /IN 0 C3225X5R1H106K250AB_p
XU4 /IN 0 C3216X7R1H105K160AE_p
R3 /RON /IN {RON}
R1 /IN /EN {REN_ADJ}
R2 /EN 0 {REN_REF}
R4 /OUT /FB {RFB_ADJ}
R5 /FB 0 {RFB_REF}
XU3 /OUT /FB C2012X7R2A223K125AE_p
V1 /IN 0 {VIN}
XU2 /SS 0 C2012X7R2A223K125AE_p
R6 /OUT 0 {RLOAD}
XU7 /OUT 0 C3216X5R0J107M160AB_p
XU5 /OUT 0 C3216X7R1H105K160AE_p
.end
